module hex7seg(input logic [3:0] hex, output logic [6:0] seg7);
    always_comb begin : sseg
        case (hex)
            4'd0:  seg7 = 7'b1000000;
            4'd1:  seg7 = 7'b0000110;
            4'd2:  seg7 = 7'b0100100;
            4'd3:  seg7 = 7'b0110000;
            4'd4:  seg7 = 7'b0011001;
            4'd5:  seg7 = 7'b0010010;
            4'd6:  seg7 = 7'b0000010;
            4'd7:  seg7 = 7'b1111000;
            4'd8:  seg7 = 7'b0000000;
            4'd9:  seg7 = 7'b0010000;
            4'd10: seg7 = 7'b0001000;
            4'd11: seg7 = 7'b0000011;
            4'd12: seg7 = 7'b1000110;
            4'd13: seg7 = 7'b0100001;
            4'd14: seg7 = 7'b0000110;
            4'd15: seg7 = 7'b0001110;
            default : seg7 = 7'b1111111;
        endcase
    end
endmodule

